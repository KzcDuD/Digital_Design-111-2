module Full_adder();